module Decoder(
    /* verilator lint_off UNUSED */
    input i_clk,
    input i_reset_n
    /* verilator lint_on UNUSED */
);


endmodule
